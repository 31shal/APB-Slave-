interface apb_intf(input clk,input reset);
  logic paddr;
  logic pwdata;
  logic psel;
  logic penable;
  logic prdata;
  logic prdata;
  logic pready;
  logic pwrite;
endinterface
